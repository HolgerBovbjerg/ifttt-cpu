mega_prog_mem_inst : mega_prog_mem PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
