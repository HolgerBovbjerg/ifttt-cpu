library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

-- 256x32 PROGRAM_MEMORY in VHDL
entity PROGRAM_MEMORY is
port(
 i_FLASH_PM_address: in std_logic_vector(7 downto 0); -- Address to read in memory 
 i_FLASH_PM_clk: in std_logic; -- clock input for FLASH_PM
 o_FLASH_PM_IR_data: out std_logic_vector(31 downto 0) -- Data output of FLASH_PM
);
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is
 
type RAM_ARRAY is array (0 to 255) of std_logic_vector (31 downto 0);


signal RAM: RAM_ARRAY :=(
-- Input in HEXADECIMAL

 	x"F0000000",x"0F000000",x"00F00000",x"000F0000",-- memory lecation 1 to 4
	x"000F0000",x"0000F000",x"0F0F0000",x"FF000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",-- memory lecation 28 to 32
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000",
	x"00000000",x"00000000",x"00000000",x"00000000"
	
	
	); 

begin
process(i_FLASH_PM_clk)
begin
 if(rising_edge(i_FLASH_PM_clk)) then
 o_FLASH_PM_IR_data <= RAM(to_integer(unsigned(i_FLASH_PM_address)));
end if;
 
end process;
 
end Behavioral;

