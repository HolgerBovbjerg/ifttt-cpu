library ieee;
use ieee.std_logic_1164.all;

package display_constants is

constant A:				std_logic_vector(7 downto 0) := x"41";
constant B:				std_logic_vector(7 downto 0) := x"42";
constant C:				std_logic_vector(7 downto 0) := x"43";
constant D:				std_logic_vector(7 downto 0) := x"44";
constant E:				std_logic_vector(7 downto 0) := x"45";
constant F:				std_logic_vector(7 downto 0) := x"46";
constant G:				std_logic_vector(7 downto 0) := x"47";
constant H:				std_logic_vector(7 downto 0) := x"48";
constant I:				std_logic_vector(7 downto 0) := x"49";
constant J:				std_logic_vector(7 downto 0) := x"4A";
constant K:				std_logic_vector(7 downto 0) := x"4B";
constant L:				std_logic_vector(7 downto 0) := x"4C";
constant M:				std_logic_vector(7 downto 0) := x"4D";
constant N:				std_logic_vector(7 downto 0) := x"4E";
constant O:				std_logic_vector(7 downto 0) := x"4F";
constant P:				std_logic_vector(7 downto 0) := x"50";
constant Q:				std_logic_vector(7 downto 0) := x"51";
constant R:				std_logic_vector(7 downto 0) := x"52";
constant S:				std_logic_vector(7 downto 0) := x"53";
constant T:				std_logic_vector(7 downto 0) := x"54";
constant U:				std_logic_vector(7 downto 0) := x"55";
constant V:				std_logic_vector(7 downto 0) := x"56";
constant W:				std_logic_vector(7 downto 0) := x"57";
constant X:				std_logic_vector(7 downto 0) := x"58";
constant Y:				std_logic_vector(7 downto 0) := x"59";
constant Z:				std_logic_vector(7 downto 0) := x"5A";
constant Zero:			std_logic_vector(7 downto 0) := x"30";
constant One:			std_logic_vector(7 downto 0) := x"31";
constant Two:			std_logic_vector(7 downto 0) := x"32";
constant Three:		std_logic_vector(7 downto 0) := x"33";
constant Four:			std_logic_vector(7 downto 0) := x"34";
constant Five:			std_logic_vector(7 downto 0) := x"35";
constant Six:			std_logic_vector(7 downto 0) := x"36";
constant Seven:		std_logic_vector(7 downto 0) := x"37";
constant Eight:		std_logic_vector(7 downto 0) := x"38";
constant Nine:			std_logic_vector(7 downto 0) := x"39";
constant Newline:		std_logic_vector(7 downto 0) := x"0A";
constant Space:		std_logic_vector(7 downto 0) := x"20";
constant Colon:		std_logic_vector(7 downto 0) := x"3A";
constant Unknown:		std_logic_vector(7 downto 0) := x"3F";

end display_constants;
package body display_constants is
end display_constants;